`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:10:13 03/29/2017 
// Design Name: 
// Module Name:    fifo_block 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fifo_top(
    output [15:0] d_rd,
    input [15:0] d_wr,
    input [7:0] a_rd,
    input [7:0] a_wr,
    input rd_en,
    input wr_en,
    input clk,
    input rst
    );



endmodule

//------------------------------------------------------
